`define CTRL_OFF  3'b000
`define CTRL_RESET_AND_SIGNAL_IF_EQUAL  3'b001
`define CTRL_COUNTDOWN_AND_SIGNAL_IF_EQUAL  3'b010
