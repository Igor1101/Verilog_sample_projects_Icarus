`define SHREG_MODE_HZ 2'b0
`define SHREG_MODE_